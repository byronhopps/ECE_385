typedef enum {UP = 0, DOWN = 1, LEFT = 2, RIGHT = 3} DIRECTION;

typedef enum {RED = 24'hFF0000, GREEN = 24'h00FF00,
    BLUE = 24'h0000FF} COLOR_24;

typedef enum {RED = 0, GREEN = 1, BLUE = 2,
    BULLET, BACKGROUND} COLOR;
