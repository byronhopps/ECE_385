module Player (
    input  logic frameClk, reset_h, clk,
    input  logic moveUp, moveDown, moveLeft, moveRight,
